`include "defines.sv"

// =============================================================================
// DCache - Phase 5: Complete Two-Level Write-Back Cache
// =============================================================================
// L1: 1KB, Direct-Mapped, LUTRAM, 16-byte lines
// - Read operations: cache enabled
// - Write hit: update L1 data, set dirty=1
// - Write miss: write-allocate (evict dirty → L2, L2 lookup → refill → write L1)
// - Eviction: if dirty, writeback to L2 (not memory)
// 
// L2: 32KB, 4-Way Set-Associative, BRAM, 16-byte lines
// - L1 miss → L2 lookup (1 cycle BRAM latency)
// - L2 hit → fill L1, return data
// - L2 miss → if victim dirty, writeback to memory; fetch from memory, fill L2+L1
// - L1 dirty eviction → UPDATE L2 entry, set L2 dirty bit
// =============================================================================

module dcache (
    input  logic        clk,
    input  logic        rst,

    // CPU Interface
    input  logic [31:0] mem_req_addr_i,
    input  logic [31:0] mem_req_wdata_i,
    input  logic        mem_req_we_i,
    input  logic [3:0]  mem_req_be_i,
    input  logic        mem_req_valid_i,

    output logic [31:0] mem_resp_data_o,
    output logic        mem_req_ready_o,
    
    // FENCE.I Cache Flush Interface
    input  logic        flush_req_i,      // Request DCache flush (all dirty lines writeback)
    output logic        flush_done_o,     // Flush operation complete

    // PTW Interface (for MMU page table walk) - Phase 1: 空实现
    input  logic [31:0] ptw_addr_i,       // PTW 请求地址
    input  logic        ptw_req_i,        // PTW 请求有效
    output logic [31:0] ptw_data_o,       // PTW 返回数据
    output logic        ptw_ack_o,        // PTW 完成应答

    // Wishbone Master Interface
    output logic [31:0] wb_adr_o,
    output logic [31:0] wb_dat_o,
    input  logic [31:0] wb_dat_i,
    output logic        wb_we_o,
    output logic [3:0]  wb_sel_o,
    output logic        wb_stb_o,
    input  logic        wb_ack_i,
    output logic        wb_cyc_o,
    input  logic        wb_rty_i,
    input  logic        wb_err_i
);

    // ========================================================================
    // L1 Cache Parameters
    // ========================================================================
    // 1KB = 64 sets × 16 bytes/line, Direct-Mapped
    localparam L1_SETS = 64;
    localparam L1_LINE_SIZE = 16;       // 16 bytes = 4 words
    localparam L1_INDEX_WIDTH = 6;      // log2(64)
    localparam L1_OFFSET_WIDTH = 4;     // log2(16)
    localparam L1_TAG_WIDTH = 22;       // 32 - 6 - 4
    localparam L1_WORD_OFFSET_WIDTH = 2;

    // ========================================================================
    // L2 Cache Parameters (Phase 4)
    // ========================================================================
    // L2_SETS can be 256 (16KB) or 512 (32KB) - other params auto-computed
    localparam L2_SETS = 256;
    localparam L2_WAYS = 4;
    localparam L2_LINE_SIZE = 16;       // 16 bytes = 4 words
    localparam L2_OFFSET_WIDTH = 4;     // log2(16) = 4
    localparam L2_INDEX_WIDTH = $clog2(L2_SETS);  // 9 for 512 sets, 8 for 256 sets
    localparam L2_TAG_WIDTH = 32 - L2_INDEX_WIDTH - L2_OFFSET_WIDTH;
    localparam L2_WORD_OFFSET_WIDTH = 2;

    // ========================================================================
    // Request Source Selection (for internal arbitration)
    // ========================================================================
    logic [31:0] current_req_addr;
    logic        current_req_valid;
    logic        current_req_we;
    logic [3:0]  current_req_be;
    logic [31:0] current_req_wdata;
    logic        current_req_is_ptw;
    
    // Priority: CPU Memory Request > PTW Request
    always_comb begin
        if (mem_req_valid_i) begin
            current_req_addr   = mem_req_addr_i;
            current_req_wdata  = mem_req_wdata_i;
            current_req_we     = mem_req_we_i;
            current_req_be     = mem_req_be_i;
            current_req_valid  = 1'b1;
            current_req_is_ptw = 1'b0;
        end else if (ptw_req_i) begin
            current_req_addr   = ptw_addr_i;
            current_req_wdata  = 32'h0;
            current_req_we     = 1'b0;      // PTW is read-only
            current_req_be     = 4'hF;      // PTW always reads full word
            current_req_valid  = 1'b1;
            current_req_is_ptw = 1'b1;
        end else begin
            current_req_addr   = 32'h0;
            current_req_wdata  = 32'h0;
            current_req_we     = 1'b0;
            current_req_be     = 4'h0;
            current_req_valid  = 1'b0;
            current_req_is_ptw = 1'b0;
        end
    end

    // ========================================================================
    // Address Breakdown
    // ========================================================================
    // L1: [31:10] Tag (22 bits) | [9:4] Index (6 bits) | [3:2] Word (2 bits) | [1:0] Byte (2 bits)
    wire [L1_TAG_WIDTH-1:0]        l1_tag   = current_req_addr[31:10];
    wire [L1_INDEX_WIDTH-1:0]      l1_index = current_req_addr[9:4];
    wire [L1_WORD_OFFSET_WIDTH-1:0] l1_word  = current_req_addr[3:2];
    
    // L2: Tag | Index | Word | Byte (widths computed from L2_SETS)
    wire [L2_TAG_WIDTH-1:0]        l2_tag   = current_req_addr[31:L2_INDEX_WIDTH+L2_OFFSET_WIDTH];
    wire [L2_INDEX_WIDTH-1:0]      l2_index = current_req_addr[L2_INDEX_WIDTH+L2_OFFSET_WIDTH-1:L2_OFFSET_WIDTH];
    wire [L2_WORD_OFFSET_WIDTH-1:0] l2_word  = current_req_addr[3:2];

    // ========================================================================
    // Address Classification
    // ========================================================================

    // Cacheable range: 0x80000000~0x807fffff (8MB)
    wire is_cacheable = (current_req_addr[31:23] == 9'b1000_0000_0);

    // ========================================================================
    // L1 Cache Storage (LUTRAM - Distributed RAM)
    // ========================================================================
    (* ram_style = "distributed" *) logic [127:0] l1_data [L1_SETS-1:0];
    (* ram_style = "distributed" *) logic [L1_TAG_WIDTH-1:0] l1_tag_array [L1_SETS-1:0];
    logic l1_valid [L1_SETS-1:0];
    logic l1_dirty [L1_SETS-1:0];  // Dirty bits for write-back

    // ========================================================================
    // L2 Cache Storage (BRAM - Block RAM)
    // ========================================================================
    // CRITICAL for BRAM inference:
    // 1. Each way needs its own array (not multi-dimensional)
    // 2. No async reset initialization (use valid bits for cold start)
    // 3. Synchronous read with output register
    
    // L2 Data arrays - one per way for BRAM inference
    (* ram_style = "block" *) logic [127:0] l2_data_way0 [L2_SETS-1:0];
    (* ram_style = "block" *) logic [127:0] l2_data_way1 [L2_SETS-1:0];
    (* ram_style = "block" *) logic [127:0] l2_data_way2 [L2_SETS-1:0];
    (* ram_style = "block" *) logic [127:0] l2_data_way3 [L2_SETS-1:0];
    
    // L2 Tag arrays - one per way for BRAM inference
    (* ram_style = "block" *) logic [L2_TAG_WIDTH-1:0] l2_tag_way0 [L2_SETS-1:0];
    (* ram_style = "block" *) logic [L2_TAG_WIDTH-1:0] l2_tag_way1 [L2_SETS-1:0];
    (* ram_style = "block" *) logic [L2_TAG_WIDTH-1:0] l2_tag_way2 [L2_SETS-1:0];
    (* ram_style = "block" *) logic [L2_TAG_WIDTH-1:0] l2_tag_way3 [L2_SETS-1:0];
    
    // Valid/Dirty bits use registers (too small for BRAM, needs async reset)
    (* ram_style = "distributed" *) logic l2_valid [L2_WAYS-1:0][L2_SETS-1:0];
    (* ram_style = "distributed" *) logic l2_dirty [L2_WAYS-1:0][L2_SETS-1:0];
    
    // LRU bits - distributed RAM or registers
    logic [2:0] l2_lru [L2_SETS-1:0];

    // ========================================================================
    // L1 Cache Lookup (Combinational - for single-cycle hit)
    // ========================================================================
    wire l1_tag_match = (l1_tag_array[l1_index] == l1_tag);
    wire l1_hit = l1_valid[l1_index] && l1_tag_match && is_cacheable;
    
    // Extract word from cache line
    logic [31:0] l1_hit_data;
    always_comb begin
        case (l1_word)
            2'b00: l1_hit_data = l1_data[l1_index][31:0];
            2'b01: l1_hit_data = l1_data[l1_index][63:32];
            2'b10: l1_hit_data = l1_data[l1_index][95:64];
            2'b11: l1_hit_data = l1_data[l1_index][127:96];
        endcase
    end

    // ========================================================================
    // L2 Cache Lookup Logic (Phase 4)
    // ========================================================================
    // L2 BRAM has 1-cycle read latency. We latch the lookup index/tag and 
    // check against BRAM outputs in next cycle.
    
    logic [L2_INDEX_WIDTH-1:0] l2_lookup_index;
    logic [L2_TAG_WIDTH-1:0]   l2_lookup_tag;
    logic [L2_WORD_OFFSET_WIDTH-1:0] l2_lookup_word;
    
    // BRAM read outputs (registered)
    logic [127:0] l2_data_read [L2_WAYS-1:0];
    logic [L2_TAG_WIDTH-1:0] l2_tag_read [L2_WAYS-1:0];
    logic l2_valid_read [L2_WAYS-1:0];
    logic l2_dirty_read [L2_WAYS-1:0];  // Phase 5: dirty bits from BRAM
    
    // L2 hit detection (combinational on registered BRAM outputs)
    logic [L2_WAYS-1:0] l2_way_hit;
    logic l2_hit;
    logic [1:0] l2_hit_way;
    logic [127:0] l2_hit_data;
    
    always_comb begin
        l2_hit = 1'b0;
        l2_hit_way = 2'b00;
        l2_hit_data = 128'h0;
        
        for (int w = 0; w < L2_WAYS; w++) begin
            l2_way_hit[w] = l2_valid_read[w] && (l2_tag_read[w] == l2_lookup_tag);
            if (l2_way_hit[w]) begin
                l2_hit = 1'b1;
                l2_hit_way = w[1:0];
                l2_hit_data = l2_data_read[w];
            end
        end
    end
    
    // Phase 5: L2 victim dirty detection (for L2 miss case)
    // Victim is selected by pseudo-LRU when we need to allocate new entry
    wire [1:0] l2_victim_way_comb = get_lru_victim(l2_lru[l2_lookup_index]);
    wire l2_victim_dirty = l2_valid_read[l2_victim_way_comb] && l2_dirty_read[l2_victim_way_comb];
    
    // Phase 5: L1 invalidation check for inclusive cache property
    // When L2 evicts a victim, must check if L1 holds that line
    // If yes, must invalidate L1 (and writeback if dirty) to maintain inclusivity
    wire [31:0] l2_victim_addr = {l2_tag_read[l2_victim_way_comb], l2_lookup_index, 4'b0000};
    wire [L1_INDEX_WIDTH-1:0] l1_victim_index = l2_victim_addr[9:4];
    wire [L1_TAG_WIDTH-1:0]   l1_victim_tag   = l2_victim_addr[31:10];
    
    // Check if L1 holds the L2 victim line
    wire l1_holds_l2_victim = l2_valid_read[l2_victim_way_comb] &&
                               l1_valid[l1_victim_index] && 
                               (l1_tag_array[l1_victim_index] == l1_victim_tag);
    wire l1_victim_needs_wb = l1_holds_l2_victim && l1_dirty[l1_victim_index];
    
    // L2 writeback data storage (latched when entering L2_WRITEBACK)
    logic [L2_TAG_WIDTH-1:0] l2_wb_tag;
    logic [127:0] l2_wb_data;
    
    // ========================================================================
    // Pseudo-LRU Functions (3-bit tree for 4-way)
    // ========================================================================
    // Tree structure:     [2]
    //                    /   \
    //                  [1]   [0]
    //                 /  \   /  \
    //              Way0 Way1 Way2 Way3
    
    function automatic logic [1:0] get_lru_victim(input logic [2:0] lru);
        if (lru[2] == 0) begin  // Go left subtree
            return lru[1] ? 2'b00 : 2'b01;
        end else begin          // Go right subtree
            return lru[0] ? 2'b10 : 2'b11;
        end
    endfunction
    
    function automatic logic [2:0] update_lru(input logic [2:0] old_lru, input logic [1:0] way);
        logic [2:0] new_lru;
        new_lru = old_lru;
        case (way)
            2'b00: begin new_lru[2] = 1'b1; new_lru[1] = 1'b1; end  // Way 0: point away
            2'b01: begin new_lru[2] = 1'b1; new_lru[1] = 1'b0; end  // Way 1: point away
            2'b10: begin new_lru[2] = 1'b0; new_lru[0] = 1'b1; end  // Way 2: point away
            2'b11: begin new_lru[2] = 1'b0; new_lru[0] = 1'b0; end  // Way 3: point away
        endcase
        return new_lru;
    endfunction


    // ========================================================================
    // FSM States
    // ========================================================================
    typedef enum logic [3:0] {
        IDLE,
        REFILL,         // Legacy: Direct L1 refill from memory (Phase 1-3)
        BYPASS_OP,      // Bypass operation (non-cacheable)
        L1_TO_L2,       // Phase 5: Write dirty L1 line to L2 (was WRITEBACK)
        L2_LOOKUP,      // Phase 4-5: Wait for L2 BRAM read (1 cycle)
        L2_REFILL,      // Phase 4-5: Fetch from memory to fill L2 (4 beats)
        L2_WRITEBACK,   // Phase 5: Write dirty L2 victim to memory (4 beats)
        L1_VICTIM_WB,   // Phase 5: Write L1 victim dirty data to L2 before L2 eviction
        FLUSH_SCAN,     // FENCE.I: Scan L1 for dirty entries
        FLUSH_L2_WB,    // FENCE.I: Write dirty L1 data to L2 (1 cycle for L2 BRAM read)
        FLUSH_WB        // FENCE.I: Writeback dirty L1 entry to memory (4 beats)
    } state_t;
    
    state_t state, next_state;

    // ========================================================================
    // Refill Logic
    // ========================================================================
    logic [1:0] refill_counter;
    logic [127:0] refill_data;

    // Latched request info (for multi-cycle operations)
    logic [31:0] latched_addr;
    logic [31:0] latched_wdata;
    logic        latched_we;
    logic [3:0]  latched_be;
    logic        latched_is_ptw;
    logic [L1_INDEX_WIDTH-1:0] latched_index;
    logic [L1_TAG_WIDTH-1:0]   latched_tag;
    logic [L1_WORD_OFFSET_WIDTH-1:0] latched_word;
    
    // Eviction address info
    logic [L1_TAG_WIDTH-1:0] old_tag;
    logic                    is_dirty_eviction;
    
    // FENCE.I Flush state
    logic [L1_INDEX_WIDTH-1:0] flush_idx;        // Current L1 set being scanned
    logic [127:0]              flush_wb_data;    // Data to writeback during flush
    logic [L1_TAG_WIDTH-1:0]   flush_wb_tag;     // Tag for flush writeback address
    logic                      flush_in_progress;// Flush operation is active
    
    // Refill address - use latched address for multi-cycle safety
    // CRITICAL: Must use latched_addr, not mem_req_addr_i, because CPU may
    // change the address during multi-cycle REFILL operation
    wire [31:0] refill_addr = {latched_addr[31:4], 4'b0000};
    
    // Writeback address - use old tag and latched index
    wire [31:0] wb_evict_addr = {old_tag, latched_index, 4'b0000};
    
    // Flush writeback address - use flush_wb_tag and flush_idx
    wire [31:0] flush_wb_addr = {flush_wb_tag, flush_idx, 4'b0000};


    // ========================================================================
    // FSM State Register
    // ========================================================================
    always_ff @(posedge clk or posedge rst) begin
        if (rst) begin
            state <= IDLE;
        end else begin
            state <= next_state;
        end
    end

    // ========================================================================
    // Request Latching
    // ========================================================================
    // Latch on:
    // 1. Cache miss (read or write)
    // 2. Write hit (for write-through operation)
    wire need_latch = current_req_valid && 
                      (!l1_hit || (l1_hit && current_req_we));
    
    always_ff @(posedge clk) begin
        if (state == IDLE && need_latch) begin
            latched_addr   <= current_req_addr;
            latched_wdata  <= current_req_wdata;
            latched_we     <= current_req_we;
            latched_be     <= current_req_be;
            latched_is_ptw <= current_req_is_ptw;
            latched_index  <= l1_index;
            latched_tag    <= l1_tag;
            latched_word   <= l1_word;
            
            // Capture victim info for potential eviction
            old_tag       <= l1_tag_array[l1_index];
            is_dirty_eviction <= l1_valid[l1_index] && l1_dirty[l1_index];
        end
    end

    // ========================================================================
    // FSM Next State Logic
    // ========================================================================
    always_comb begin
        next_state = state;
        
        case (state)
            IDLE: begin
                // FENCE.I flush request has priority over normal operations
                if (flush_req_i) begin
                    next_state = FLUSH_SCAN;
                end else if (current_req_valid) begin
                    if (is_cacheable) begin
                        if (l1_hit) begin
                            if (current_req_we) begin
                                // Write hit: Update L1 immediately (done in IDLE), stay in IDLE
                                // Single-cycle write using combinational signals
                                next_state = IDLE; 
                            end else begin
                                // Read hit: Return data immediately
                                next_state = IDLE;
                            end
                        end else begin
                            // L1 Miss (Read or Write)
                            // Only write dirty L1 data to L2 on eviction
                            if (l1_valid[l1_index] && l1_dirty[l1_index]) begin
                                next_state = L1_TO_L2; // Write dirty L1 line to L2
                            end else begin
                                next_state = L2_LOOKUP;  // Clean or invalid, check L2 directly
                            end
                        end
                    end else begin
                        // Non-cacheable access -> Bypass
                        next_state = BYPASS_OP;
                    end
                end
            end
            
            FLUSH_SCAN: begin
                // Scan L1 for dirty entries
                // Check if current flush_idx is dirty
                if (l1_valid[flush_idx] && l1_dirty[flush_idx]) begin
                    // Dirty entry found - first update L2, then writeback to memory
                    // L2 BRAM read is initiated on this transition (see l2_bram_rd_en logic)
                    next_state = FLUSH_L2_WB;
                end else begin
                    // Not dirty, advance to next set or finish
                    if (flush_idx == L1_SETS - 1) begin
                        // All sets scanned, flush complete
                        next_state = IDLE;
                    end
                    // else: stay in FLUSH_SCAN, flush_idx will increment
                end
            end
            
            FLUSH_L2_WB: begin
                // Wait 1 cycle for L2 BRAM read, then write L1 data to L2 and proceed to FLUSH_WB
                // L2 write happens in this state (see l2_bram_wr_en logic)
                next_state = FLUSH_WB;
            end
            
            FLUSH_WB: begin
                // Writeback dirty L1 entry to memory (4 beats)
                if (wb_ack_i && refill_counter == 2'b11) begin
                    // Writeback complete
                    if (flush_idx == L1_SETS - 1) begin
                        // All sets scanned, flush complete
                        next_state = IDLE;
                    end else begin
                        // Continue scanning
                        next_state = FLUSH_SCAN;
                    end
                end
            end
            
            L2_LOOKUP: begin
                // Wait 1 cycle for L2 BRAM read, then check hit/miss
                if (l2_hit) begin
                    // L2 hit: Fill L1 from L2, complete immediately
                    next_state = IDLE;
                end else begin
                    // L2 miss: Need to evict victim and refill
                    // Phase 5: First check if L1 has dirty data for L2 victim
                    if (l1_victim_needs_wb) begin
                        // L1 has dirty version of L2 victim - must writeback to L2 first
                        next_state = L1_VICTIM_WB;
                    end else if (l2_victim_dirty) begin
                        // L2 victim is dirty, writeback to memory
                        next_state = L2_WRITEBACK;
                    end else begin
                        // Victim is clean (or only L1 holds clean copy), proceed to refill
                        next_state = L2_REFILL;
                    end
                end
            end
            
            L2_REFILL: begin
                // Fetching from memory to fill L2 (4 beats)
                if (wb_ack_i && refill_counter == 2'b11) begin
                    // L2 refill complete, also fill L1, return to IDLE
                    next_state = IDLE;
                end
            end
            
            REFILL: begin
                // Phase 3 legacy path (direct L1 refill from memory)
                // This is still used for some scen arios
                if (wb_ack_i && refill_counter == 2'b11) begin
                    next_state = IDLE;
                end
            end
            
            BYPASS_OP: begin
                if (wb_ack_i) begin
                    next_state = IDLE;
                end
            end
            
            L1_TO_L2: begin
                // Phase 5: Single cycle write of L1 dirty line to L2
                // L2 always contains L1 (inclusive), so this is an UPDATE
                next_state = L2_LOOKUP;
            end
            
            L2_WRITEBACK: begin
                // Phase 5: Write dirty L2 victim to memory (4 beats)
                if (wb_ack_i && refill_counter == 2'b11) begin
                    // L2 writeback done, now do actual refill
                    next_state = L2_REFILL;
                end
            end
            
            L1_VICTIM_WB: begin
                // Phase 5: Single cycle write of L1 victim dirty data to L2 victim
                // This updates L2 victim with L1's dirty data before L2 eviction
                // After this, L2 victim is dirty and must be written back to memory
                next_state = L2_WRITEBACK;
            end
            
            default: next_state = IDLE;
        endcase
    end

    // ========================================================================
    // Refill Counter
    // ========================================================================
    always_ff @(posedge clk or posedge rst) begin
        if (rst) begin
            refill_counter <= 2'b00;
        end else if (state != REFILL && state != L2_REFILL && state != L2_WRITEBACK && state != FLUSH_WB) begin
            refill_counter <= 2'b00;
        end else if ((state == REFILL || state == L2_REFILL || state == L2_WRITEBACK || state == FLUSH_WB) && wb_ack_i) begin
            refill_counter <= refill_counter + 2'b01;
        end
    end
    
    // ========================================================================
    // FENCE.I Flush Index Counter and Data Latching
    // ========================================================================
    always_ff @(posedge clk or posedge rst) begin
        if (rst) begin
            flush_idx <= '0;
            flush_in_progress <= 1'b0;
            flush_wb_data <= 128'h0;
            flush_wb_tag <= '0;
        end else begin
            // Entering FLUSH_SCAN from IDLE
            if (state == IDLE && next_state == FLUSH_SCAN) begin
                flush_idx <= '0;
                flush_in_progress <= 1'b1;
            end
            // In FLUSH_SCAN, advancing to next set if current is clean
            else if (state == FLUSH_SCAN && next_state == FLUSH_SCAN) begin
                flush_idx <= flush_idx + 1'b1;
            end
            // Entering FLUSH_L2_WB - latch data and tag for L2 update and memory writeback
            else if (state == FLUSH_SCAN && next_state == FLUSH_L2_WB) begin
                flush_wb_data <= l1_data[flush_idx];
                flush_wb_tag  <= l1_tag_array[flush_idx];
            end
            // After FLUSH_WB completes, advance to next set (in FLUSH_SCAN)
            else if (state == FLUSH_WB && next_state == FLUSH_SCAN) begin
                flush_idx <= flush_idx + 1'b1;
            end
            // Flush complete - return to IDLE
            else if ((state == FLUSH_SCAN || state == FLUSH_WB || state == FLUSH_L2_WB) && next_state == IDLE) begin
                flush_in_progress <= 1'b0;
            end
        end
    end
    
    // Flush done output - asserted for one cycle when flush completes
    assign flush_done_o = flush_in_progress && (state == FLUSH_SCAN || state == FLUSH_WB) && next_state == IDLE;

    // ========================================================================
    // Refill Data Accumulation
    // ========================================================================
    always_ff @(posedge clk) begin
        if ((state == REFILL || state == L2_REFILL) && wb_ack_i) begin
            case (refill_counter)
                2'b00: refill_data[31:0]   <= wb_dat_i;
                2'b01: refill_data[63:32]  <= wb_dat_i;
                2'b10: refill_data[95:64]  <= wb_dat_i;
                2'b11: refill_data[127:96] <= wb_dat_i;
            endcase
        end
    end
    
    // ========================================================================
    // L2 BRAM Read Logic (Phase 4-5)
    // ========================================================================
    // Read from L2 BRAM when:
    // 1. Entering L2_LOOKUP: read new address to check hit/miss
    // 2. Entering L1_TO_L2: read evicted address to find target way
    // Results are available next cycle.
    
    // Compute evicted address L2 index for BRAM read
    // CRITICAL: When transitioning IDLE→L1_TO_L2, old_tag/latched_index are being latched
    // on the SAME clock edge, so we must use LIVE signals here (not latched).
    wire [L1_TAG_WIDTH-1:0] evict_tag_live = l1_tag_array[l1_index];
    wire [L2_INDEX_WIDTH-1:0] evict_l2_idx = {evict_tag_live[L2_INDEX_WIDTH-L1_INDEX_WIDTH-1:0], l1_index};
    
    always_ff @(posedge clk) begin
        if (state == IDLE && next_state == L2_LOOKUP) begin
            // Latch lookup parameters for new address
            l2_lookup_index <= l2_index;
            l2_lookup_tag   <= l2_tag;
            l2_lookup_word  <= l2_word;
        end else if (state == L1_TO_L2 && next_state == L2_LOOKUP) begin
            // After L1_TO_L2, latch lookup parameters for the NEW address
            l2_lookup_index <= l2_index;
            l2_lookup_tag   <= l2_tag;
            l2_lookup_word  <= l2_word;
        end
    end
    
    // ========================================================================
    // L2 BRAM Read Logic - Unified Address Port
    // ========================================================================
    // CRITICAL for BRAM inference: Use a SINGLE registered address for reads.
    // All read conditions feed into this address register.
    
    logic [L2_INDEX_WIDTH-1:0] l2_bram_rd_addr;
    logic l2_bram_rd_en;
    
    // Compute flush address L2 index (similar to evict_l2_idx)
    // flush_l2_addr = {flush_wb_tag, flush_idx, 4'b0000} → L2_index = addr[12:4]
    // CRITICAL: Use LIVE signals from L1 (not latched) since latch happens on same edge
    wire [L1_TAG_WIDTH-1:0] flush_tag_live = l1_tag_array[flush_idx];
    wire [L2_INDEX_WIDTH-1:0] flush_l2_idx = {flush_tag_live[L2_INDEX_WIDTH-L1_INDEX_WIDTH-1:0], flush_idx};
    wire [L2_TAG_WIDTH-1:0]   flush_l2_tag = {flush_tag_live[L1_TAG_WIDTH-1:L2_INDEX_WIDTH-L1_INDEX_WIDTH]};
    
    // Compute the read address based on state transitions
    always_comb begin
        l2_bram_rd_addr = l2_index; // default
        l2_bram_rd_en = 1'b0;
        
        if (state == IDLE && next_state == L2_LOOKUP) begin
            l2_bram_rd_addr = l2_index;
            l2_bram_rd_en = 1'b1;
        end else if (state == IDLE && next_state == L1_TO_L2) begin
            l2_bram_rd_addr = evict_l2_idx;
            l2_bram_rd_en = 1'b1;
        end else if (state == L1_TO_L2 && next_state == L2_LOOKUP) begin
            l2_bram_rd_addr = l2_index;
            l2_bram_rd_en = 1'b1;
        end else if (state == FLUSH_SCAN && next_state == FLUSH_L2_WB) begin
            // Read L2 to find which way holds the flush line
            l2_bram_rd_addr = flush_l2_idx;
            l2_bram_rd_en = 1'b1;
        end
    end
    
    // BRAM Read: Single address port, synchronous read
    always_ff @(posedge clk) begin
        if (l2_bram_rd_en) begin
            l2_data_read[0]  <= l2_data_way0[l2_bram_rd_addr];
            l2_data_read[1]  <= l2_data_way1[l2_bram_rd_addr];
            l2_data_read[2]  <= l2_data_way2[l2_bram_rd_addr];
            l2_data_read[3]  <= l2_data_way3[l2_bram_rd_addr];
            
            l2_tag_read[0]   <= l2_tag_way0[l2_bram_rd_addr];
            l2_tag_read[1]   <= l2_tag_way1[l2_bram_rd_addr];
            l2_tag_read[2]   <= l2_tag_way2[l2_bram_rd_addr];
            l2_tag_read[3]   <= l2_tag_way3[l2_bram_rd_addr];
            
            l2_valid_read[0] <= l2_valid[0][l2_bram_rd_addr];
            l2_valid_read[1] <= l2_valid[1][l2_bram_rd_addr];
            l2_valid_read[2] <= l2_valid[2][l2_bram_rd_addr];
            l2_valid_read[3] <= l2_valid[3][l2_bram_rd_addr];
            
            l2_dirty_read[0] <= l2_dirty[0][l2_bram_rd_addr];
            l2_dirty_read[1] <= l2_dirty[1][l2_bram_rd_addr];
            l2_dirty_read[2] <= l2_dirty[2][l2_bram_rd_addr];
            l2_dirty_read[3] <= l2_dirty[3][l2_bram_rd_addr];
        end
    end
    
    // Phase 5: Latch L2 victim data when entering L2_WRITEBACK
    always_ff @(posedge clk) begin
        if (state == L2_LOOKUP && next_state == L2_WRITEBACK) begin
            // Latch victim way's tag and data for memory writeback (L2 already dirty)
            l2_wb_tag  <= l2_tag_read[l2_victim_way_comb];
            l2_wb_data <= l2_data_read[l2_victim_way_comb];
        end else if (state == L1_VICTIM_WB && next_state == L2_WRITEBACK) begin
            // Coming from L1_VICTIM_WB: we just wrote L1 data to L2, writeback that
            // Tag is still the L2 victim's original tag
            l2_wb_tag  <= l2_tag_read[l2_victim_way_comb];
            l2_wb_data <= l1_victim_data_latched;  // Use REGISTERED data (latched when entering L1_VICTIM_WB)
        end
    end

    // ========================================================================
    // L1 Cache Update (on refill complete OR write-through)
    // ========================================================================
    
    // Compute new cache line for write-through (apply byte-enable mask)
    // NOTE: Use LIVE request signals (not latched) for immediate cache update
    logic [127:0] write_through_line;
    logic [31:0]  write_through_word;
    
    always_comb begin
        // Apply byte-enable to create the new word
        // Use l1_hit_data (from current address) and current request data
        write_through_word = l1_hit_data;  // Start with current cache data
        if (mem_req_be_i[0]) write_through_word[7:0]   = mem_req_wdata_i[7:0];
        if (mem_req_be_i[1]) write_through_word[15:8]  = mem_req_wdata_i[15:8];
        if (mem_req_be_i[2]) write_through_word[23:16] = mem_req_wdata_i[23:16];
        if (mem_req_be_i[3]) write_through_word[31:24] = mem_req_wdata_i[31:24];
        
        // Insert the modified word into the cache line
        // Use l1_index (current address), not latched_index
        write_through_line = l1_data[l1_index];
        case (l1_word)
            2'b00: write_through_line[31:0]   = write_through_word;
            2'b01: write_through_line[63:32]  = write_through_word;
            2'b10: write_through_line[95:64]  = write_through_word;
            2'b11: write_through_line[127:96] = write_through_word;
        endcase
    end
    
    // Refill data with write-allocate merge
    logic [127:0] refill_line_merged;
    logic [31:0]  refill_word_merged;
    logic [127:0] refill_line_full;  // Complete refill line
    
    always_comb begin
        // First, construct the COMPLETE refill line (including last beat)
        refill_line_full = {wb_dat_i, refill_data[95:0]};
        
        // Extract the target word from the complete line
        case (latched_word)
            2'b00: refill_word_merged = refill_line_full[31:0];
            2'b01: refill_word_merged = refill_line_full[63:32];
            2'b10: refill_word_merged = refill_line_full[95:64];
            2'b11: refill_word_merged = refill_line_full[127:96];
        endcase
        
        // Apply byte-enable mask for write-allocate
        if (latched_we) begin
             if (latched_be[0]) refill_word_merged[7:0]   = latched_wdata[7:0];
             if (latched_be[1]) refill_word_merged[15:8]  = latched_wdata[15:8];
             if (latched_be[2]) refill_word_merged[23:16] = latched_wdata[23:16];
             if (latched_be[3]) refill_word_merged[31:24] = latched_wdata[31:24];
        end
        
        // Construct the final merged line
        refill_line_merged = refill_line_full;
        if (latched_we) begin
             case (latched_word)
                 2'b00: refill_line_merged[31:0]   = refill_word_merged;
                 2'b01: refill_line_merged[63:32]  = refill_word_merged;
                 2'b10: refill_line_merged[95:64]  = refill_word_merged;
                 2'b11: refill_line_merged[127:96] = refill_word_merged;
             endcase
        end
    end
    
    // L2 hit write-allocate merge logic
    // This computes the merged line when an L2 hit occurs for a write request
    logic [127:0] l2_hit_line_merged;
    logic [31:0]  l2_hit_word_merged;
    
    always_comb begin
        // Extract the target word from L2 hit data
        case (latched_word)
            2'b00: l2_hit_word_merged = l2_hit_data[31:0];
            2'b01: l2_hit_word_merged = l2_hit_data[63:32];
            2'b10: l2_hit_word_merged = l2_hit_data[95:64];
            2'b11: l2_hit_word_merged = l2_hit_data[127:96];
        endcase
        
        // Apply byte-enable mask for write-allocate
        if (latched_be[0]) l2_hit_word_merged[7:0]   = latched_wdata[7:0];
        if (latched_be[1]) l2_hit_word_merged[15:8]  = latched_wdata[15:8];
        if (latched_be[2]) l2_hit_word_merged[23:16] = latched_wdata[23:16];
        if (latched_be[3]) l2_hit_word_merged[31:24] = latched_wdata[31:24];
        
        // Construct the merged line
        l2_hit_line_merged = l2_hit_data;
        case (latched_word)
            2'b00: l2_hit_line_merged[31:0]   = l2_hit_word_merged;
            2'b01: l2_hit_line_merged[63:32]  = l2_hit_word_merged;
            2'b10: l2_hit_line_merged[95:64]  = l2_hit_word_merged;
            2'b11: l2_hit_line_merged[127:96] = l2_hit_word_merged;
        endcase
    end
    
    integer i, j;
    always_ff @(posedge clk or posedge rst) begin
        if (rst) begin
            // Reset unpacked arrays with loop
            for (i = 0; i < L1_SETS; i = i + 1) begin
                l1_valid[i] <= 1'b0;
                l1_dirty[i] <= 1'b0;
            end
        end else if (state == L2_LOOKUP && l2_hit) begin
            // L2 Hit: Fill L1 from L2
            // For WRITES: Also apply write data and set dirty
            if (latched_we) begin
                // Write hit: Use pre-computed merged line (computed in always_comb below)
                l1_data[latched_index]      <= l2_hit_line_merged;
                l1_dirty[latched_index]     <= 1'b1;  // Dirty because we modified it
            end else begin
                // Read hit: Just fill L1 with L2 data
                l1_data[latched_index]      <= l2_hit_data;
                l1_dirty[latched_index]     <= 1'b0;  // Clean from L2
            end
            l1_tag_array[latched_index] <= latched_tag;
            l1_valid[latched_index]     <= 1'b1;
            
        end else if (state == L2_REFILL && wb_ack_i && refill_counter == 2'b11) begin
            // L2 Refill complete - Fill L1 from refilled data
            // Also handle write-allocate if needed
            if (latched_we) begin
                l1_data[latched_index]  <= refill_line_merged;
                l1_dirty[latched_index] <= 1'b1;  // Dirty because we modified it
            end else begin
                l1_data[latched_index]  <= {wb_dat_i, refill_data[95:0]};
                l1_dirty[latched_index] <= 1'b0;  // Clean (fresh from memory)
            end
            l1_tag_array[latched_index] <= latched_tag;
            l1_valid[latched_index]     <= 1'b1;
            
            // Phase 5: CRITICAL - Also invalidate L1 entry for L2 victim if present
            // This must be done here, not in a separate else-if branch!
            // Only invalidate if:
            // 1. L1 held the L2 victim line (l1_holds_l2_victim_latched)
            // 2. The victim index is different from the index we just filled
            //    (otherwise we'd invalidate the line we just wrote)
            if (l1_holds_l2_victim_latched && l1_victim_index_latched != latched_index) begin
                l1_valid[l1_victim_index_latched] <= 1'b0;
            end
            
        end else if (state == REFILL && wb_ack_i && refill_counter == 2'b11) begin
            // Legacy REFILL path (Phase 3 compatibility)
            // Refill complete - write cache line
            // If Write-Allocate (latched_we=1), we write the MERGED line and set DIRTY
            if (latched_we) begin
                l1_data[latched_index]  <= refill_line_merged;
                l1_dirty[latched_index] <= 1'b1;  // Dirty because we modified it
            end else begin
                l1_data[latched_index]  <= {wb_dat_i, refill_data[95:0]};
                l1_dirty[latched_index] <= 1'b0;  // Clean (fresh from memory)
            end
            l1_tag_array[latched_index] <= latched_tag;
            l1_valid[latched_index]     <= 1'b1;
            
        end else if (state == IDLE && current_req_valid && l1_hit && current_req_we && !current_req_is_ptw) begin
            // Write Hit: update L1 cache line immediately (CPU only, PTW is read-only)
            // Single-cycle operation using combinational signals
            l1_data[l1_index] <= write_through_line;
            l1_dirty[l1_index] <= 1'b1; // Mark as dirty
            
        end else if (state == L1_VICTIM_WB) begin
            // Phase 5: L1 victim writeback - invalidate L1 entry
            l1_valid[l1_victim_index] <= 1'b0;
            
        end else if (state == FLUSH_WB && wb_ack_i && refill_counter == 2'b11) begin
            // FENCE.I: Flush writeback complete - mark L1 entry as clean
            // Keep L1 valid - subsequent accesses can still hit L1.
            // L1/L2 consistency is now maintained by always writing L1 to L2 on eviction.
            l1_dirty[flush_idx] <= 1'b0;
        end
    end
    
    // ========================================================================
    // L2 Cache Update Logic (Phase 5)
    // ========================================================================
    // L2 is updated on:
    // 1. L2_REFILL completion (memory fetch) - dirty=0
    // 2. L2 hit (LRU update only)
    // 3. L1_TO_L2 (dirty L1 writeback) - dirty=1
    
    logic [1:0] l2_victim_way;
    
    // Evicted L1 line's L2 address (computed from old_tag + latched_index)
    wire [31:0] evicted_addr = {old_tag, latched_index, 4'b0000};
    wire [L2_TAG_WIDTH-1:0]   evicted_l2_tag   = evicted_addr[31:L2_INDEX_WIDTH+L2_OFFSET_WIDTH];
    wire [L2_INDEX_WIDTH-1:0] evicted_l2_index = evicted_addr[L2_INDEX_WIDTH+L2_OFFSET_WIDTH-1:L2_OFFSET_WIDTH];
    
    // L2 way that holds the evicted L1 line (for L1_TO_L2 update)
    // Since L2 is inclusive, the evicted line MUST be in L2
    // We use the l2_lookup results which were read when entering L1_TO_L2
    logic [1:0] l1_to_l2_target_way;
    logic l1_to_l2_found;
    
    // Combinational logic to find which L2 way has the evicted line
    always_comb begin
        l1_to_l2_found = 1'b0;
        l1_to_l2_target_way = 2'b00;
        for (int w = 0; w < L2_WAYS; w++) begin
            if (l2_valid_read[w] && (l2_tag_read[w] == evicted_l2_tag)) begin
                l1_to_l2_found = 1'b1;
                l1_to_l2_target_way = w[1:0];
            end
        end
    end
    
    // L1 data to write to L2 (captured when entering L1_TO_L2)
    logic [127:0] l1_evicted_data;
    always_ff @(posedge clk) begin
        if (state == IDLE && next_state == L1_TO_L2) begin
            l1_evicted_data <= l1_data[l1_index];
        end
    end
    
    // FLUSH_L2_WB: Find which L2 way holds the flush line
    // Similar to l1_to_l2_found but uses flush_l2_tag (latched as flush_wb_tag)
    logic [1:0] flush_l2_target_way;
    logic flush_l2_way_found;
    wire [L2_TAG_WIDTH-1:0] flush_l2_tag_latched = flush_wb_tag[L1_TAG_WIDTH-1:L2_INDEX_WIDTH-L1_INDEX_WIDTH];
    wire [L2_INDEX_WIDTH-1:0] flush_l2_idx_latched = {flush_wb_tag[L2_INDEX_WIDTH-L1_INDEX_WIDTH-1:0], flush_idx};
    
    always_comb begin
        flush_l2_way_found = 1'b0;
        flush_l2_target_way = 2'b00;
        for (int w = 0; w < L2_WAYS; w++) begin
            if (l2_valid_read[w] && (l2_tag_read[w] == flush_l2_tag_latched)) begin
                flush_l2_way_found = 1'b1;
                flush_l2_target_way = w[1:0];
            end
        end
    end
    
    // L2 valid/dirty reset logic (separate from BRAM writes)
    always_ff @(posedge clk or posedge rst) begin
        if (rst) begin
            for (i = 0; i < L2_SETS; i = i + 1) begin
                l2_lru[i] <= 3'b000;
                for (j = 0; j < L2_WAYS; j = j + 1) begin
                    l2_valid[j][i] <= 1'b0;
                    l2_dirty[j][i] <= 1'b0;
                end
            end
        end else if (state == L1_TO_L2) begin
            // Phase 5: Update valid/dirty/LRU for L1->L2 writeback
            if (l1_to_l2_found) begin
                // Only set L2 dirty if L1 was dirty (is_dirty_eviction is latched on L1 miss)
                // If L1 was clean, L2 should remain clean to avoid spurious memory writebacks
                l2_dirty[l1_to_l2_target_way][evicted_l2_index] <= is_dirty_eviction;
                l2_lru[evicted_l2_index] <= update_lru(l2_lru[evicted_l2_index], l1_to_l2_target_way);
            end
        end else if (state == L2_LOOKUP && l2_hit) begin
            // L2 Hit: Update LRU
            l2_lru[l2_lookup_index] <= update_lru(l2_lru[l2_lookup_index], l2_hit_way);
        end else if (state == L1_VICTIM_WB) begin
            // Phase 5: Update L2 dirty bit (L1 valid invalidation moved to L1 Update block)
            l2_dirty[l2_victim_way_comb][l2_lookup_index] <= 1'b1;
        end else if (state == L2_REFILL && wb_ack_i && refill_counter == 2'b11) begin
            // L2 Refill complete: Update valid/dirty/LRU
            // Note: L1 valid invalidation moved to L1 Update block
            l2_victim_way = get_lru_victim(l2_lru[l2_lookup_index]);
            l2_valid[l2_victim_way][l2_lookup_index] <= 1'b1;
            l2_dirty[l2_victim_way][l2_lookup_index] <= 1'b0;
            l2_lru[l2_lookup_index] <= update_lru(l2_lru[l2_lookup_index], l2_victim_way);
        end else if (state == FLUSH_L2_WB && flush_l2_way_found) begin
            // FLUSH_L2_WB: Update L2 with dirty L1 data, set dirty=0 (will write to memory next)
            l2_dirty[flush_l2_target_way][flush_l2_idx_latched] <= 1'b0;
            l2_lru[flush_l2_idx_latched] <= update_lru(l2_lru[flush_l2_idx_latched], flush_l2_target_way);
        end
    end
    
    // ========================================================================
    // L2 BRAM Write Logic - Unified Interface
    // ========================================================================
    // CRITICAL for BRAM inference: Use unified write address/data/enable signals
    // to ensure single-port write behavior.
    
    logic l2_bram_wr_en;
    logic [L2_INDEX_WIDTH-1:0] l2_bram_wr_addr;
    logic [127:0] l2_bram_wr_data;
    logic [L2_TAG_WIDTH-1:0] l2_bram_wr_tag;
    logic [1:0] l2_bram_wr_way;
    logic l2_bram_wr_tag_en;  // Only write tag on refill, not on updates
    
    // Compute write signals based on state
    always_comb begin
        l2_bram_wr_en = 1'b0;
        l2_bram_wr_addr = l2_lookup_index;
        l2_bram_wr_data = 128'h0;
        l2_bram_wr_tag = l2_lookup_tag;
        l2_bram_wr_way = 2'b00;
        l2_bram_wr_tag_en = 1'b0;
        
        if (state == L1_TO_L2 && l1_to_l2_found) begin
            // Write dirty L1 data to L2 (update existing entry)
            l2_bram_wr_en = 1'b1;
            l2_bram_wr_addr = evicted_l2_index;
            l2_bram_wr_data = l1_evicted_data;
            l2_bram_wr_way = l1_to_l2_target_way;
            l2_bram_wr_tag_en = 1'b0;  // Don't update tag (already correct)
        end else if (state == L1_VICTIM_WB) begin
            // Write L1 victim dirty data to L2 victim way
            // CRITICAL: Use latched data instead of dynamic l1_data[l1_victim_index]
            l2_bram_wr_en = 1'b1;
            l2_bram_wr_addr = l2_lookup_index;
            l2_bram_wr_data = l1_victim_data_latched;  // Use REGISTERED data
            l2_bram_wr_way = l2_victim_way_comb;
            l2_bram_wr_tag_en = 1'b0;  // Don't update tag
        end else if (state == L2_REFILL && wb_ack_i && refill_counter == 2'b11) begin
            // L2 refill complete - write new line
            // CRITICAL FIX: For write-allocate, use refill_line_merged (with write data merged)
            // to ensure L1 and L2 have consistent data. Previously used raw refill data which
            // would contain undefined values for uninitialized memory addresses.
            l2_bram_wr_en = 1'b1;
            l2_bram_wr_addr = l2_lookup_index;
            l2_bram_wr_data = latched_we ? refill_line_merged : {wb_dat_i, refill_data[95:0]};
            l2_bram_wr_way = get_lru_victim(l2_lru[l2_lookup_index]);
            l2_bram_wr_tag = l2_lookup_tag;
            l2_bram_wr_tag_en = 1'b1;  // Update tag
        end else if (state == FLUSH_L2_WB && flush_l2_way_found) begin
            // FLUSH_L2_WB: Update L2 with dirty L1 data before writing to memory
            l2_bram_wr_en = 1'b1;
            l2_bram_wr_addr = flush_l2_idx_latched;
            l2_bram_wr_data = flush_wb_data;
            l2_bram_wr_way = flush_l2_target_way;
            l2_bram_wr_tag_en = 1'b0;  // Don't update tag (already correct)
        end
    end
    
    // BRAM Write: Data arrays - Single always block with case statement
    // Write on: L1_TO_L2, L1_VICTIM_WB, L2_REFILL
    always_ff @(posedge clk) begin
        if (l2_bram_wr_en) begin
            case (l2_bram_wr_way)
                2'b00: l2_data_way0[l2_bram_wr_addr] <= l2_bram_wr_data;
                2'b01: l2_data_way1[l2_bram_wr_addr] <= l2_bram_wr_data;
                2'b10: l2_data_way2[l2_bram_wr_addr] <= l2_bram_wr_data;
                2'b11: l2_data_way3[l2_bram_wr_addr] <= l2_bram_wr_data;
            endcase
        end
    end
    
    // BRAM Write: Tag arrays - Separate always block, only on L2_REFILL
    always_ff @(posedge clk) begin
        if (l2_bram_wr_en && l2_bram_wr_tag_en) begin
            case (l2_bram_wr_way)
                2'b00: l2_tag_way0[l2_bram_wr_addr] <= l2_bram_wr_tag;
                2'b01: l2_tag_way1[l2_bram_wr_addr] <= l2_bram_wr_tag;
                2'b10: l2_tag_way2[l2_bram_wr_addr] <= l2_bram_wr_tag;
                2'b11: l2_tag_way3[l2_bram_wr_addr] <= l2_bram_wr_tag;
            endcase
        end
    end
    
    // Phase 5: Latch L1 victim info when entering various states
    logic l1_holds_l2_victim_latched;
    logic [L1_INDEX_WIDTH-1:0] l1_victim_index_latched;
    logic [127:0] l1_victim_data_latched;  // NEW: Latch L1 victim data for BRAM write
    
    always_ff @(posedge clk) begin
        if (state == L2_LOOKUP && next_state == L2_REFILL) begin
            l1_holds_l2_victim_latched <= l1_holds_l2_victim;
            l1_victim_index_latched <= l1_victim_index;
        end else if (state == L2_LOOKUP && next_state == L2_WRITEBACK) begin
            // Also latch when going to L2_WRITEBACK (will eventually go to L2_REFILL)
            l1_holds_l2_victim_latched <= l1_holds_l2_victim;
            l1_victim_index_latched <= l1_victim_index;
        end else if (state == L2_LOOKUP && next_state == L1_VICTIM_WB) begin
            // Latch L1 victim data BEFORE entering L1_VICTIM_WB state
            // This is CRITICAL for BRAM inference - eliminates dynamic combinational access
            l1_holds_l2_victim_latched <= l1_holds_l2_victim;
            l1_victim_index_latched <= l1_victim_index;
            l1_victim_data_latched <= l1_data[l1_victim_index];  // Latch the data
        end
    end

    // ========================================================================
    // Wishbone Interface
    // ========================================================================
    always_comb begin
        wb_we_o  = 1'b0;
        wb_sel_o = 4'b1111;
        wb_stb_o = 1'b0;
        wb_cyc_o = 1'b0;
        wb_adr_o = 32'h0;
        wb_dat_o = 32'h0;
        
        case (state)
            REFILL: begin
                wb_adr_o = refill_addr + {28'b0, refill_counter, 2'b00};
                wb_we_o  = 1'b0;
                wb_sel_o = 4'b1111;
                wb_stb_o = 1'b1;
                wb_cyc_o = 1'b1;
            end
           
            L2_REFILL: begin
                // Fetch from memory to fill L2 (Phase 4)
                wb_adr_o = refill_addr + {28'b0, refill_counter, 2'b00};
                wb_we_o  = 1'b0;
                wb_sel_o = 4'b1111;
                wb_stb_o = 1'b1;
                wb_cyc_o = 1'b1;
            end
            
            BYPASS_OP: begin
                wb_adr_o = latched_addr;
                wb_dat_o = latched_wdata;
                wb_we_o  = latched_we;
                wb_sel_o = latched_be;
                wb_stb_o = 1'b1;
                wb_cyc_o = 1'b1;
            end
            
            L2_WRITEBACK: begin
                // Phase 5: Write dirty L2 victim line back to memory
                // L2 victim address constructed from l2_lookup (tag + index)
                wb_adr_o = {l2_wb_tag, l2_lookup_index, 4'b0000} + {28'b0, refill_counter, 2'b00};
                wb_we_o  = 1'b1;
                wb_sel_o = 4'b1111;
                wb_stb_o = 1'b1;
                wb_cyc_o = 1'b1;
                
                // Select word to write from L2 victim data
                case (refill_counter)
                    2'b00: wb_dat_o = l2_wb_data[31:0];
                    2'b01: wb_dat_o = l2_wb_data[63:32];
                    2'b10: wb_dat_o = l2_wb_data[95:64];
                    2'b11: wb_dat_o = l2_wb_data[127:96];
                endcase
            end
            
            FLUSH_WB: begin
                // FENCE.I: Write dirty L1 entry to memory (4 beats)
                wb_adr_o = flush_wb_addr + {28'b0, refill_counter, 2'b00};
                wb_we_o  = 1'b1;
                wb_sel_o = 4'b1111;
                wb_stb_o = 1'b1;
                wb_cyc_o = 1'b1;
                
                // Select word to write from flushed L1 data
                case (refill_counter)
                    2'b00: wb_dat_o = flush_wb_data[31:0];
                    2'b01: wb_dat_o = flush_wb_data[63:32];
                    2'b10: wb_dat_o = flush_wb_data[95:64];
                    2'b11: wb_dat_o = flush_wb_data[127:96];
                endcase
            end
            
            default: begin
                // IDLE, L1_TO_L2, L2_LOOKUP, FLUSH_SCAN - no wishbone activity
            end
        endcase
    end

    // ========================================================================
    // Response Data Selection
    // ========================================================================
    // CRITICAL: refill_data has been updated in previous cycles via non-blocking
    // assignment, so it's valid to read. For word 3 on beat 3, use wb_dat_i directly.
    logic [31:0] refill_word;
    always_comb begin
        case (latched_word)
            2'b00: refill_word = refill_data[31:0];     // Word 0 was loaded at beat 0
            2'b01: refill_word = refill_data[63:32];    // Word 1 was loaded at beat 1
            2'b10: refill_word = refill_data[95:64];    // Word 2 was loaded at beat 2
            2'b11: refill_word = wb_dat_i;              // Word 3 is current beat (beat 3)
        endcase
    end

    // ========================================================================
    // Output Mux
    // ========================================================================
    // Internal combinational signals for PTW response
    logic [31:0] ptw_data_comb;
    logic        ptw_ack_comb;
    
    always_comb begin
        mem_resp_data_o = 32'h0;
        mem_req_ready_o = 1'b0;
        ptw_data_comb   = 32'h0;
        ptw_ack_comb    = 1'b0;
        
        if (state == IDLE && current_req_valid && l1_hit && !current_req_we) begin
            // L1 read hit - immediate response
            if (current_req_is_ptw) begin
                ptw_data_comb = l1_hit_data;
                ptw_ack_comb  = 1'b1;
            end else begin
                mem_resp_data_o = l1_hit_data;
                mem_req_ready_o = 1'b1;
            end
        end else if (state == IDLE && current_req_valid && l1_hit && current_req_we) begin
            // Write hit - immediate completion (L1 updated in FF)
            // CPU only, PTW doesn't write
            mem_resp_data_o = 32'h0;
            mem_req_ready_o = 1'b1;
        end else if (state == L2_LOOKUP && l2_hit) begin
            // L2 hit - return requested word from L2
            logic [31:0] l2_hit_word;
            case (l2_lookup_word)
                2'b00: l2_hit_word = l2_hit_data[31:0];
                2'b01: l2_hit_word = l2_hit_data[63:32];
                2'b10: l2_hit_word = l2_hit_data[95:64];
                2'b11: l2_hit_word = l2_hit_data[127:96];
            endcase
            if (latched_is_ptw) begin
                ptw_data_comb = l2_hit_word;
                ptw_ack_comb  = 1'b1;
            end else begin
                mem_resp_data_o = l2_hit_word;
                mem_req_ready_o = 1'b1;
            end
        end else if (state == L2_REFILL && wb_ack_i && refill_counter == 2'b11) begin
            // L2 Refill complete - return requested word
            if (latched_is_ptw) begin
                ptw_data_comb = refill_word;
                ptw_ack_comb  = 1'b1;
            end else begin
                mem_resp_data_o = refill_word;
                mem_req_ready_o = 1'b1;
            end
        end else if (state == REFILL && wb_ack_i && refill_counter == 2'b11) begin
            // Legacy REFILL complete - return requested word
            if (latched_is_ptw) begin
                ptw_data_comb = refill_word;
                ptw_ack_comb  = 1'b1;
            end else begin
                mem_resp_data_o = refill_word;
                mem_req_ready_o = 1'b1;
            end
        end else if (state == BYPASS_OP && wb_ack_i) begin
            // Bypass operation complete
            if (latched_is_ptw) begin
                ptw_data_comb = wb_dat_i;
                ptw_ack_comb  = 1'b1;
            end else begin
                mem_resp_data_o = wb_dat_i;
                mem_req_ready_o = 1'b1;
            end
        end
    end
    
    // ========================================================================
    // PTW Response Delay Register (1 cycle)
    // ========================================================================
    // This delay is CRITICAL for ptw_arbiter and MMU timing:
    // - Allows ptw_arbiter state machine to update before ack arrives
    // - Allows MMU to enter LEVEL1_WAIT/LEVEL2_WAIT before seeing ack
    always_ff @(posedge clk or posedge rst) begin
        if (rst) begin
            ptw_data_o <= 32'h0;
            ptw_ack_o  <= 1'b0;
        end else begin
            ptw_data_o <= ptw_data_comb;
            ptw_ack_o  <= ptw_ack_comb;
        end
    end

endmodule
